LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE work.aux_package.all;
USE ieee.numeric_std.ALL;
--USE ieee.std_logic_ARITH.all;
use ieee.std_logic_unsigned.all;
-------------------------------------
ENTITY ALU IS
  generic (
		n : positive := 8 ; -- A,B length
		m : positive := 5 ; -- OPC length
		k : positive := 2   -- STATUS length
	);
  PORT (    cin : IN STD_LOGIC;
			A,B : in std_logic_vector(n-1 downto 0);
			OPC : in std_logic_vector(m-1 downto 0);

		----------------------------------------
			RES : out std_logic_vector(2*n-1 downto 0); -- Result(HI,LO)
			STATUS : out std_logic_vector(k-1 downto 0));
END ALU;
------------- complete the top Architecture code --------------
ARCHITECTURE struct OF ALU IS


	SIGNAL ACC : std_logic_vector(2*n-1 DOWNTO 0):=(others=> '0'); -- for the BarrelShfter
	--SIGNAL Result:std_logic_vector(2*n-1 downto 0);
	--adder:
	Signal sel:std_logic_vector(1 downto 0);
	Signal adderRes:std_logic_vector(n-1 downto 0);
	signal adderCout:std_logic;
BEGIN

--AddSub:Adder generic map (n) port map (cin,A,B,sel,adderCout,adderRes);

PROCESS (OPC,A,B,cin)
variable Along,Blong,Result:std_logic_vector(2*n-1 downto 0);
variable AccVar,tmp:std_logic_vector(2*n DOWNTO 0);


	BEGIN
	
	Along:=(others=> '0');
	Blong:=(others=> '0');
	Along(n-1 downto 0) := A;
	Blong(n-1 downto 0) := B;
	
	Result := ( others => '0');
	STATUS <= "00";

	  	case OPC(4 downto 0) is
		  when "00001" =>   Result := Along+Blong;
							--sel <= "00";
							--Result(n downto 0) := adderCout & adderRes;
							
		  when "00010" =>   Result := Along-Blong;
							--sel <= "10";
							--Result(n downto 0) := adderCout & adderRes;
		  when "00011" =>   Result := Along+Blong+cin;
		  					--sel <= "01";
							--Result(n downto 0) := adderCout & adderRes;
		  when "00100" =>   Result := std_logic_vector(unsigned(A)*unsigned(B));
		  
		  when "00101" =>   AccVar := ( others => '0');
							AccVar(2*n-1 downto 0) := std_logic_vector(unsigned(A)*unsigned(B));							
							
							if (AccVar + ACC) < 2**(2*n) - 1  then -- check if Acc makes CARRY and zeroes him
							AccVar := AccVar + ACC;
							ACC <=AccVar(2*n-1 DOWNTO 0);
							Result := AccVar(2*n-1 DOWNTO 0);

							else
							STATUS(0) <= '1';
							tmp := (AccVar + ACC) -2**(2*n);
							Result := tmp(2*n-1 DOWNTO 0);
							ACC<= (others=> '0');
							end if;						
							
							
		  when "00110" =>   ACC <= (others=>'0'); --acc Resultet
		  when "00111" => if A<B then
							Result := Blong; --max
							else Result := Along;
							end if;
							
		  when "01000" => if A<B then
				Result := Along; --min
				else Result := Blong;
				end if;
			when "01001" => --and
						Result(n-1 downto 0) := A and B;				
			when "01010" => -- or
						Result(n-1 downto 0) := A or B;
			when "01011" =>	--xor	
						Result(n-1 downto 0) := A xor B;			
		   when others => Result := (others=> '1'); --not for me 
		end case;
		
		if Result = 0 then 
			STATUS(1) <= '1';
		end if;
				
		RES <= Result; -- we used an internal signal Result
	END PROCESS;
	
	
	
	
	
	

END struct;

--configure list -delta collapse